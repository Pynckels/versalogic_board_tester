* 2N3906 PNP Transistor SPICE Model
.model 2N3906 PNP (IS=1.89f BF=200 NF=1.0 VAF=20 IKF=0.05 XTB=1.5 BR=3 NR=1.0 VAR=10 IKR=0.03 RC=1.0 CJE=6p VJE=0.75 MJE=0.333 CJC=4p VJC=0.75 MJC=0.333 TF=0.8n TR=40n)
