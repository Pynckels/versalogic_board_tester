.SUBCKT BS250P D G S
Cgs  G S 20.1E-12
Cgd1 G 4 57.1E-12
Cgd2 D 4 5E-12
M1 D G S S MOST1
M2 4 G D S MOST2
D1 D S Dbody
.ENDS

.MODEL MOST1 PMOS(LEVEL=3 VTO=-2.3 W=7.6m L=2u KP=10.33u RD=4.014 RS=20m)
.MODEL MOST2 PMOS(VTO=2.43 W=7.6m L=2u KP=10.33u RS=20m)
.MODEL Dbody D(CJO=53.22E-12 VJ=0.5392 M=0.3583 IS=75.32E-15 N=1.016 RS=1.245 TT=86.56n BV=45 IBV=10u
