* 2N3904 NPN Transistor SPICE Model
.model 2N3904 NPN (IS=6.734f BF=416.4 NF=1.0 VAF=74.03 IKF=0.284 XTB=1.5 BR=3.162 NR=1.0 VAR=12.63 IKR=0.03 RC=1.0 CJE=4.3p VJE=0.75 MJE=0.333 CJC=2.2p VJC=0.75 MJC=0.333 TF=0.984n TR=35.05n)
