
* VO1400 SPICE MODEL
*							LED ANODE
*							| LED Cathode
*							| |  Pin 4 SSR contact
*							| |  |  Pin 3 SSR contact
*							| |  |  |
*							| |  |  |

.SUBCKT VO1400              A C  S1 S2

* Simplified model of the input LED and its forward voltage
D1 A V_LED_IN D_IDEAL
R_ON V_LED_IN C 1k
V_IN V_LED_IN 0 DC 0

* Voltage-controlled switch for the output
S1 S1 S2 V_IN C SW_MODEL

* Passive components for robustness
R_LEAK S1 S2 10G
C_PARASITIC S1 S2 1p
.ENDS

.model D_IDEAL D(Is=1p)
.model SW_MODEL VSWITCH(Ron=1 Roff=10G Voff=2.0 Von=3.5)
