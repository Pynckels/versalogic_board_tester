* G3VM-41AY1-compatible opto-MOSFET relay model
* Pins: 1=A (Anode), 2=K (Cathode), 3=D (Drain), 4=S (Source)

.subckt G3VM-41AY1 A K D S

* LED diode model (approx. VF = 1.27V @10mA)
DLED A K D_LED
RLED A K 2        ; Rs = 2Ω series resistance

.model D_LED D(IS=8e-16 N=1.7 RS=0)

* RC delay to simulate switching time (2.8ms ON, 0.3ms OFF)
Rdelay A nctrl 1k
Cdelay nctrl K 1u

* Voltage-controlled switch as output FET
* Controlled by voltage across LED via RC node
S1 D S nctrl K SMOS

.model SMOS VSWITCH(Ron=0.09 Roff=1Meg Vt=1 Vh=0.1)

.ends G3VM-41AY1
