* ADG417 SPICE Macro-model (Fixed for ngspice compatibility)
* Compatible with KiCad 9 + ngspice

* Force ngspice to accept behavioral expressions
.option numdgt=7
.option ngbehavior=ps

* Pinout:
*      1  = S1
*      2  = NC
*      3  = GND
*      4  = VDD
*      5  = RESET/VL
*      6  = IN1
*      7  = VSS
*      8  = D1

* Switch Models
.MODEL VON     SW(VT=0.8 VH=0.1 RON=0.001     ROFF=1.8E8)
.MODEL VEN     SW(VT=0.8 VH=0.1 RON=1.073E5   ROFF=1.1621E5)
.MODEL VRESET  SW(VT=0.8 VH=0.1 RON=2.7E6     ROFF=1K)
.MODEL DCLAMP  D(IS=1E-15 IBV=1E-13)

.SUBCKT ADG417 1 3 4 5 6 7 8

* RESET/VL
S30 5 187 5 3 VRESET
C80 187 3 5.5E-11

* IDD/ISS
I1 4 3 1E-10
I2 7 3 1E-10

* ESD PROTECTION DIODES
D11 7 8 DCLAMP
D12 8 4 DCLAMP
D13 7 1 DCLAMP
D14 1 4 DCLAMP

* OFF ISOLATION
C11 1 8 3.2E-13

* CHARGE INJECTION
C12 8 140 2.3E-12
C13 1 140 2.3E-12

* CD/CS OFF AND BANDWIDTH
C14 1 3 1E-12
C15 8 3 1E-12

* ON RESISTANCE SWITCHING LOGIC
Ech155 1555 3 VALUE = { IF(ABS(V(1)) > ABS(V(184)), V(1), V(8)) }
R155 1555 3 1G
R11 137 8 0.001

S111 136 141 1141 3 VON
Ech111 1141 3 VALUE = { IF(V(1555) < -11.9339, 5, 0) }
Ech11 141 3 VALUE = { IF(V(1555) < -11.9339, 0.193250257331202 * (V(1555) + 11.9339) + 23.7255, 0) }

S112 136 146 1146 3 VON
Ech112 1146 3 VALUE = { IF(V(1555) >= -11.9339 && V(1555) <= 13.8208, 5, 0) }
Ech12 146 3 VALUE = { IF(V(1555) >= -11.9339 && V(1555) <= 13.8208, ((23.7255 - 15.1961) / ((-11.9339 - 2.77905599210194)^2)) * (V(1555) - 2.77905599210194)^2 + 15.1961, 0) }

S113 136 144 1144 3 VON
Ech113 1144 3 VALUE = { IF(V(1555) > 13.8208, 5, 0) }
Ech13 144 3 VALUE = { IF(V(1555) > 13.8208, -0.219543147208122 * (V(1555) - 13.8208) + 20, 0) }

RIN1 136 3 1G
EOUT1 137 181 VALUE = { V(136,3) * 0.000999 }
FCOPY1 3 180 VSENSE1 1
RSENSOR1 180 3 1K
VSENSE1 181 184 DC 0

* TON / TOFF / BBM
S11 182 184 140 3 VON
S12 143 138 143 3 VEN
Ech14 143 3 VALUE = { 2.9 + 2.1 * tanh((2.4-V(6))/0.1) }
* Fixed EV1 definition to avoid poly source ambiguity
EV1 140 3 VALUE = { V(138,3) }
C16 138 3 1E-12

* VOLTAGE SUPPLY REQUIREMENTS
S13 1 182 185 3 VON
S14 142 185 142 3 VON
Ech15 142 3 VALUE = { IF((V(7) <= -0.5 && V(7) >= -16.5) && (V(4) <= 16.5 && V(4) >= 5), 5, 0.01) }
S15 139 185 139 3 VON
Ech16 139 3 VALUE = { IF(V(7) >= -0.5 && V(4) <= 16.5 && V(4) >= 5, 5, 0.01) }

.ENDS ADG417
